module bcd_comparator();

endmodule